module ReservationStation (
    input   clk, rst_n, enable
);
    
endmodule