module lsq #(
    parameters
) (
    ports
);
    
endmodule